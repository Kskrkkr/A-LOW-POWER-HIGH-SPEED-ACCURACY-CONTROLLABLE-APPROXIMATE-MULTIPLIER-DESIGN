`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.10.2025 17:35:24
// Design Name: 
// Module Name: testbench64
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench64;
reg [63:0]r;
reg [5:0]sel;
wire y;

mux_64a testbench(.a(r[63:0]),.sel(sel[5:0]),.y(y));

initial
begin

sel=6'b000000; r=64'b0000000000000000000000000000000000000000000000000000000000000001;#10
sel=6'b000101; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b001001; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b000001; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b000001; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b110001; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b000001; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b000111; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b011001; r=64'b0000000000000000000000000000000000000000000000000000000000000101;#10
sel=6'b111111; r=64'b1111111111111111111111111111111111111111111111111111111111111111;#10
$stop;

end
endmodule
